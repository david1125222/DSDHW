module barrel_shifter(in, shift, out);
input  [7:0] in;
input  [2:0] shift;
output [7:0] out;

/*Write your code here*/
assign output = (shift==3'h0) ? 

/*End of code*/
endmodule